
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0] in1;
    logic [7:0] in2;
    logic   add_sub;
    logic [8:0] out;
    //--------------------------------------------------------------------------

endinterface

